module top_module ( input a, input b, output out );
    mod_a instance_mod_a(a, b, out);
endmodule

